module ddk

// 	//todo safe ordered concurrent map
