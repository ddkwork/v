module demo

// 	//todo safe ordered concurrent map
