module ddk
