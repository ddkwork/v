module demo
